typedef enum logic [4:0] {
    SMState0,
    SMState1,
    SMState2,
    SMState3,
    SMState4,
    SMState5,
    SMReset,
    SimResetting,
    SMResetComplete,
    SMIdle
} SimState /*verilator public*/; 
