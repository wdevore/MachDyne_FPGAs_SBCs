// `define FIRMWARE "../binaries/firmware.hex"
`define FIRMWARE "/media/RAMDisk/firmware.hex"

