typedef enum logic [4:0] {
    SMState0,
    SMState1,
    SMState2,
    SMState3,
    SMState4,
    SMState5,
    SMState6,
    SMState7,
    SMReset,
    SimResetting,
    SMResetComplete,
    SMIdle   // 11
} SimState /*verilator public*/; 
