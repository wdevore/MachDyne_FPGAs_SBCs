    SMEnableInterrupts_S1,  // 4
    SMEnableInterrupts_S2,  // 5
    SMEnableInterrupts_S3,  // 6

    SMEnableInterrupts_S4,  // 7
    SMEnableInterrupts_S5,  // 8
    SMEnableInterrupts_S6,  // 9
    SMEnableInterrupts_S7,  // 10
    SMEnableInterrupts_S8,  // 11
    SMEnableInterrupts_S9,  // 12
    SMEnableInterrupts_S10,  // 13
    SMEnableInterrupts_S11,  // 14
    SMEnableInterrupts_S12,  // 15
    SMEnableInterrupts_S13,  // 16
    SMEnableInterrupts_S14,  // 17
    SMEnableInterrupts_S15,  // 18
    SMEnableInterrupts_S16,  // 19
