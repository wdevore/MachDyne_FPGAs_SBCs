    SM_S1,   // 4
    SM_S2,   // 5
    SM_S3,
    
    SM_S4,

    SM_S5,
    SM_S6,
    SM_S7,

    SM_S8,
    SM_S9,
    SM_S10,
    SM_S11,

    SM_S12,

    // SMStop // 20
