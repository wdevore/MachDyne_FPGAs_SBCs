typedef enum logic [2:0] {
    UAReset0,
    UAReset1,
    UAResetComplete
} UARTState; 
