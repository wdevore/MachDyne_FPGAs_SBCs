typedef enum logic [2:0] {
    SMReset0,
    SMReset1,
    SMResetComplete
} SimState; 
