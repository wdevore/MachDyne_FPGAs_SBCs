`define FIRMWARE "/media/RAMDisk/firmware.hex"

`define SYSCLK 50_000_000
`define SDRAM_CLK_FREQ (`SYSCLK / 1_000_000)

