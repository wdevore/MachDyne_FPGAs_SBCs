    SM_S1,   // 4
    SM_S2,   // 5
    SM_S3,
    SM_S4,
    SM_S5,

    // SMStop // 20
