typedef enum logic [4:0] {
    SMReset,
    SMResetComplete,
    SMIdle,
    Vector2,
    Vector3
} SimState /*verilator public*/; 
