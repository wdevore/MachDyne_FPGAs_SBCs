`define FIRMWARE "../../binaries/firmware.hex"

