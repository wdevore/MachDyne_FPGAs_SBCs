typedef enum logic [4:0] {
    SMReset,
    SMResetComplete,
    SMIdle
} SimState /*verilator public*/; 
