    SMClientRejection_S1,   // 4
    SMClientRejection_S2,   // 5
    SMClientRejection_S3,
    SMClientRejection_S4,

    SMClientRejection_S5,
    SMClientRejection_S6,
    SMClientRejection_S7,
    SMClientRejection_S8,

    SMClientRejection_S9, 
    SMClientRejection_S10,
    SMClientRejection_S11,

    SMClientRejection_S12,
    SMClientRejection_S13,
    SMClientRejection_S14,
    SMClientRejection_S15,

    SMClientRejection_S16,
    SMClientRejection_S17,
    SMClientRejection_S18,  // 21

    // SMStop // 20
