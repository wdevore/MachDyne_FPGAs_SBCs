// Defines specific to the Schoko.
// Most of these are deprecated in favor of simply copying 
// everything needed from sysctl_pico.v

`define FPGA_ECP5
`define OSC48
`define SYSCLK50
`define VCLK25
`define EN_SDRAM
`define EN_BSRAM32
`define EN_UART0

`define FIRMWARE_PATH "../MiniSchoko/gas/sdram/"