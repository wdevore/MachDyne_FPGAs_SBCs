typedef enum logic [5:0] {
    RAMState0,
    RAMState1,
    RAMState2,
    SDReset,
    SDResetting,
    SDIdle
} SDRAMState;

